module hello; endmodule
