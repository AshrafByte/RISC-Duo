`default_nettype none
import types_pkg::*;
import types_pkg::*;
