`default_nettype none

module newmod; endmodule
