`default_nettype none
import types_pkg::*;

module testmod; endmodule
