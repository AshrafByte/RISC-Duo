`default_nettype none
import types_pkg::*;

